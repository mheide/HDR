library ieee;
use ieee.std_logic_1164.all;

entity test_exposure_control is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity test_exposure_control;

architecture RTL of test_exposure_control is
	
begin

end architecture RTL;
